thermal grid 1
R12 1 2 1
R23 2 3 1
R45 4 5 1
R56 5 6 1
R78 7 8 1
R89 8 9 1
R14 1 4 1
R47 4 7 1
R25 2 5 1
R58 5 8 1
R36 3 6 1
R69 6 9 1
VAMB 9 0 300
I1  0 1 1
I2  0 2 1
I3  0 3 1
I4  0 4 1
I5  0 5 1
I6  0 6 1
I7  0 7 1
I8  0 8 1
I9  0 9 1
.print dc v(*)
.op
.end